`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/15/2020 07:26:12 PM
// Design Name: 
// Module Name: Learning_random
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Learning_random(
    input [3:0] a,b,
    output [4:0] y
    );
    
    assign y=a+b;
    
    
endmodule
