`include "uvm_macros.svh"
import uvm_pkg::*;

class transaction extends uvm_sequence_item;
rand bit[3:0] a;
rand bit [7:0] b;
function new(input string inst="TRANS");
super.new(inst);
endfunction
`uvm_object_utils_begin(transaction)
`uvm_field_int(a,UVM_DEFAULT)
`uvm_field_int(b,UVM_DEFAULT)
`uvm_object_utils_end
endclass

class producer extends uvm_component;
`uvm_component_utils(producer)
transaction t;
integer i;

uvm_blocking_put_port #(transaction) send;

function new(input string inst="PROD", uvm_component c);
super.new(inst,c);
send=new("PUT",this);
endfunction
virtual function void build_phase(uvm_phase phase);
super.build_phase(phase);
t=transaction::type_id::create("TRANS",this);
endfunction

virtual task run_phase(uvm_phase phase);
phase.raise_objection(phase);
for(i=0;i<10;i++) begin
#40;
t.randomize();
`uvm_info("PROD","Data sent",UVM_NONE);
t.print(uvm_default_line_printer);
send.put(t);
end
phase.drop_objection(phase);
endtask
endclass

class consumer extends uvm_component;
`uvm_component_utils(consumer)
transaction data;
integer i;

uvm_blocking_get_port #(transaction) recv;

function new(input string inst="CONS", uvm_component c);
super.new(inst,c);
recv=new("GET",this);
endfunction

virtual function void build_phase(uvm_phase phase);
super.build_phase(phase);
data=transaction::type_id::create("TRANS",this);
endfunction

virtual task run_phase(uvm_phase phase);
phase.raise_objection(phase);
for(i=0;i<10;i++) begin
#40;
recv.get(data);
`uvm_info("CONS",$sformatf("Data received : %0d",data),UVM_NONE);
data.print(uvm_default_line_printer);
end
phase.drop_objection(phase);
endtask
endclass

class env extends uvm_env;
`uvm_component_utils(env)

producer p; 
consumer c;
uvm_tlm_fifo #(transaction) fifo;
function new(input string inst="ENV", uvm_component c);
super.new(inst,c);
endfunction

virtual function void build_phase(uvm_phase phase);
super.build_phase(phase);
p=producer::type_id::create("PROD",this);
c=consumer::type_id::create("CONS",this);
fifo=new("FIFO",this,1);
endfunction

virtual function void connect_phase(uvm_phase phase);
super.connect_phase(phase);
p.send.connect(fifo.put_export);
c.recv.connect(fifo.get_export);
endfunction

virtual task run_phase(uvm_phase phase);
forever begin
#40;
if(fifo.is_full())
begin
`uvm_info("ENV","Fifo is full",UVM_NONE);
end
else begin
`uvm_info("ENV","Fifo is not full",UVM_NONE);
end
end
endtask
endclass

class test extends uvm_test;
`uvm_component_utils(test)
env e;
function new(string inst="TEST",uvm_component c);
super.new(inst,c);
endfunction
virtual function void build_phase(uvm_phase phase);
super.build_phase(phase);
e=env::type_id::create("ENV",this);
endfunction

endclass

module tb;
test t;
initial begin
t=new("TEST",null);
run_test();
end
endmodule